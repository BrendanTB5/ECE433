`timescale 1ns / 100ps
//Brendan Mulholland CM1832
//ECE343 HW2 Problem 7
//9/22/19
//This is the Test Bench for Detect 1001

module hw2p7BNMTest;

	// Inputs
	
      
endmodule

